module geofence ( clk,reset,X,Y,valid,is_inside);
input clk;
input reset;
input [9:0] X;
input [9:0] Y;
output valid;
output is_inside;
//reg valid;
//reg is_inside;
reg [3:0] hello_world ;
reg[4:0] ll;
reg[4:0] hh;



endmodule
